package Parameters;
//Parameters for encoding and decoding needs to stay the same
parameter SEARCH_BUFFER_DEPTH = 8;
parameter SEARCH_BUFFER_WIDTH = 7;
parameter SEARCH_BUFFER_SIZE = SEARCH_BUFFER_DEPTH*SEARCH_BUFFER_WIDTH; 
parameter LOOKAHEAD_BUFFER_LENGTH = 6;
parameter SYMBOL_LENGTH = 8;

endpackage